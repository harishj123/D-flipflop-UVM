//interface
interface dff_interface(input logic clk);
  logic rst;
  logic din;
  logic dout;
endinterface
